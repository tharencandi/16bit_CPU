module lab5_part3(clk,out,clr);

output[15:0] out;
input clk,clr;
wire[25:0] Q;
reg Enable;

fiftyMHz_counter inst_count1(.clk(clk),.Q(Q),.clr(clr));

always @(posedge clk) begin
	if (Q == 26'd0)
		Enable <= 1'b1;
		
	else
		Enable <= 1'b0;
end

sixteenb_counter inst_count2(.Enable(Enable), .clk(clk), .clr(clr), .Q(out));

endmodule