module program_counter(clk, rst, bus, select, enable);
	
	input bus, 



	

	
