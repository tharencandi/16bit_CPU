module output_sig(state, out);

input [3:0] state;
output reg out;

always @(state) begin
	case (state)
	4'b0100 : begin out = 1'b1; end
	4'b1000 : begin out = 1'b1; end
	default : begin out = 1'b0; end
	
	endcase
	end
	
endmodule